/***** SDRAM COMMANDS *****/
`define CMD_COMMAND_INHIBIT 	 0
`define CMD_NOP			    	 1
`define CMD_ACTIVE			 	 2
`define CMD_READ					 3
`define CMD_WRITE					 4
`define CMD_BURST_TERMINATE 	 5
`define CMD_PRECHARGE		 	 6
`define CMD_AUTO_REFRESH	 	 7
`define CMD_LOAD_MODE_REGISTER 8