/**** ACTIONS ON ADDRESS AND BANK BUSES ****/
`define CLEAR_A_B		  0 
`define SET_A_10		  1
`define CLEAR_A		  2
`define MODE_REG_SETUP 3
`define ASSIGN_WR_PTR  4
`define ASSIGN_RD_PTR  5